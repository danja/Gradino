**************************************************************
*  Electronic circuit simulation file                        *
*                                                            *
**************************************************************

* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
* SUBCKT TL071   1 2 3 4 5

.INCLUDE bits.mod  

* Low pass

Rsrc 0 1 1K
C1 1 2 1UF
R1 2 3 10K
X1 0 3 20 21 4 TL071

R2 3 4 47K
C2 3 4 4.7n

R3 10 8 10K

* extra
R8 4 10 10K
* C4 10 0 560p
C4 10 12 100n
R10 12 0 5.6K

* High Pass
C3 1 5 5.6n
* C3 1 5 10n
R4 5 6 10K
X2 0 6 20 21 7 TL071
R5 6 7 47K

* extra
* C5 7 11 100n
R9 7 11 0
* C5 7 11 1n

* mix
R6 11 8 10K
R7 8 9 10K
X3 0 8 20 21 9 TL071

Vcc 20 0 15
Vee 21 0 -15

Vsrc  1  0   dc 0   ac 1 

* Vsrc	1	0	SIN(0V .1VPEAK 1KHZ)
* .TRAN 	10US 1000US


.control
* .AC DEC 10000 1u 1Meg 
AC DEC 10 10 1MEGHZ
plot vdb(9)
.endc
.END

